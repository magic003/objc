module runtime

pub type Bool = bool

pub const yes = Bool(true)

pub const no = Bool(false)
