module runtime

type Id = C.objc_object
