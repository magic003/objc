module objc

// A type that represents a Boolean value in Objective-C.
pub type Bool = bool

// yes as true.
pub const yes = Bool(true)

// no as false.
pub const no = Bool(false)
