module main

fn main() {
	app := TrayApp.new()
	app.init()
	app.run()
}
